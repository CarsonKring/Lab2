module stimulus;